`include "defines.v"


module sha1(

    input wire clk,
    input wire rst
    );

endmodule
