`include "defines.v"


module sha1(

    input wire clk,
    // input wire rst,
    input wire[`Sha1In] sha1_i,         // 从外设读取的数据
    output wire[`Sha1Out] sha1_o        // 读、写外设的地址
    );

    reg [`Sha1Pad] sha_pad;

    reg[31:0] W[80:0];
    reg[31:0] A[80:0];
    reg[31:0] B[80:0];
    reg[31:0] C[80:0];
    reg[31:0] D[80:0];
    reg[31:0] E[80:0];
    reg[31:0] TEMP[80:0];
    
wire[31:0] w0;
wire[31:0] w1;
wire[31:0] w2;
wire[31:0] w3;
wire[31:0] w4;
wire[31:0] w5;
wire[31:0] w6;
wire[31:0] w7;
wire[31:0] w8;
wire[31:0] w9;
wire[31:0] w10;
wire[31:0] w11;
wire[31:0] w12;
wire[31:0] w13;
wire[31:0] w14;
wire[31:0] w15;
wire[31:0] w16;
wire[31:0] w17;
wire[31:0] w18;
wire[31:0] w19;
wire[31:0] w20;
wire[31:0] w21;
wire[31:0] w22;
wire[31:0] w23;
wire[31:0] w24;
wire[31:0] w25;
wire[31:0] w26;
wire[31:0] w27;
wire[31:0] w28;
wire[31:0] w29;
wire[31:0] w30;
wire[31:0] w31;
wire[31:0] w32;
wire[31:0] w33;
wire[31:0] w34;
wire[31:0] w35;
wire[31:0] w36;
wire[31:0] w37;
wire[31:0] w38;
wire[31:0] w39;
wire[31:0] w40;
wire[31:0] w41;
wire[31:0] w42;
wire[31:0] w43;
wire[31:0] w44;
wire[31:0] w45;
wire[31:0] w46;
wire[31:0] w47;
wire[31:0] w48;
wire[31:0] w49;
wire[31:0] w50;
wire[31:0] w51;
wire[31:0] w52;
wire[31:0] w53;
wire[31:0] w54;
wire[31:0] w55;
wire[31:0] w56;
wire[31:0] w57;
wire[31:0] w58;
wire[31:0] w59;
wire[31:0] w60;
wire[31:0] w61;
wire[31:0] w62;
wire[31:0] w63;
wire[31:0] w64;
wire[31:0] w65;
wire[31:0] w66;
wire[31:0] w67;
wire[31:0] w68;
wire[31:0] w69;
wire[31:0] w70;
wire[31:0] w71;
wire[31:0] w72;
wire[31:0] w73;
wire[31:0] w74;
wire[31:0] w75;
wire[31:0] w76;
wire[31:0] w77;
wire[31:0] w78;
wire[31:0] w79;
wire[31:0] w80;
wire[31:0] a0;
wire[31:0] a1;
wire[31:0] a2;
wire[31:0] a3;
wire[31:0] a4;
wire[31:0] a5;
wire[31:0] a6;
wire[31:0] a7;
wire[31:0] a8;
wire[31:0] a9;
wire[31:0] a10;
wire[31:0] a11;
wire[31:0] a12;
wire[31:0] a13;
wire[31:0] a14;
wire[31:0] a15;
wire[31:0] a16;
wire[31:0] a17;
wire[31:0] a18;
wire[31:0] a19;
wire[31:0] a20;
wire[31:0] a21;
wire[31:0] a22;
wire[31:0] a23;
wire[31:0] a24;
wire[31:0] a25;
wire[31:0] a26;
wire[31:0] a27;
wire[31:0] a28;
wire[31:0] a29;
wire[31:0] a30;
wire[31:0] a31;
wire[31:0] a32;
wire[31:0] a33;
wire[31:0] a34;
wire[31:0] a35;
wire[31:0] a36;
wire[31:0] a37;
wire[31:0] a38;
wire[31:0] a39;
wire[31:0] a40;
wire[31:0] a41;
wire[31:0] a42;
wire[31:0] a43;
wire[31:0] a44;
wire[31:0] a45;
wire[31:0] a46;
wire[31:0] a47;
wire[31:0] a48;
wire[31:0] a49;
wire[31:0] a50;
wire[31:0] a51;
wire[31:0] a52;
wire[31:0] a53;
wire[31:0] a54;
wire[31:0] a55;
wire[31:0] a56;
wire[31:0] a57;
wire[31:0] a58;
wire[31:0] a59;
wire[31:0] a60;
wire[31:0] a61;
wire[31:0] a62;
wire[31:0] a63;
wire[31:0] a64;
wire[31:0] a65;
wire[31:0] a66;
wire[31:0] a67;
wire[31:0] a68;
wire[31:0] a69;
wire[31:0] a70;
wire[31:0] a71;
wire[31:0] a72;
wire[31:0] a73;
wire[31:0] a74;
wire[31:0] a75;
wire[31:0] a76;
wire[31:0] a77;
wire[31:0] a78;
wire[31:0] a79;
wire[31:0] a80;
wire[31:0] b0;
wire[31:0] b1;
wire[31:0] b2;
wire[31:0] b3;
wire[31:0] b4;
wire[31:0] b5;
wire[31:0] b6;
wire[31:0] b7;
wire[31:0] b8;
wire[31:0] b9;
wire[31:0] b10;
wire[31:0] b11;
wire[31:0] b12;
wire[31:0] b13;
wire[31:0] b14;
wire[31:0] b15;
wire[31:0] b16;
wire[31:0] b17;
wire[31:0] b18;
wire[31:0] b19;
wire[31:0] b20;
wire[31:0] b21;
wire[31:0] b22;
wire[31:0] b23;
wire[31:0] b24;
wire[31:0] b25;
wire[31:0] b26;
wire[31:0] b27;
wire[31:0] b28;
wire[31:0] b29;
wire[31:0] b30;
wire[31:0] b31;
wire[31:0] b32;
wire[31:0] b33;
wire[31:0] b34;
wire[31:0] b35;
wire[31:0] b36;
wire[31:0] b37;
wire[31:0] b38;
wire[31:0] b39;
wire[31:0] b40;
wire[31:0] b41;
wire[31:0] b42;
wire[31:0] b43;
wire[31:0] b44;
wire[31:0] b45;
wire[31:0] b46;
wire[31:0] b47;
wire[31:0] b48;
wire[31:0] b49;
wire[31:0] b50;
wire[31:0] b51;
wire[31:0] b52;
wire[31:0] b53;
wire[31:0] b54;
wire[31:0] b55;
wire[31:0] b56;
wire[31:0] b57;
wire[31:0] b58;
wire[31:0] b59;
wire[31:0] b60;
wire[31:0] b61;
wire[31:0] b62;
wire[31:0] b63;
wire[31:0] b64;
wire[31:0] b65;
wire[31:0] b66;
wire[31:0] b67;
wire[31:0] b68;
wire[31:0] b69;
wire[31:0] b70;
wire[31:0] b71;
wire[31:0] b72;
wire[31:0] b73;
wire[31:0] b74;
wire[31:0] b75;
wire[31:0] b76;
wire[31:0] b77;
wire[31:0] b78;
wire[31:0] b79;
wire[31:0] b80;
wire[31:0] c0;
wire[31:0] c1;
wire[31:0] c2;
wire[31:0] c3;
wire[31:0] c4;
wire[31:0] c5;
wire[31:0] c6;
wire[31:0] c7;
wire[31:0] c8;
wire[31:0] c9;
wire[31:0] c10;
wire[31:0] c11;
wire[31:0] c12;
wire[31:0] c13;
wire[31:0] c14;
wire[31:0] c15;
wire[31:0] c16;
wire[31:0] c17;
wire[31:0] c18;
wire[31:0] c19;
wire[31:0] c20;
wire[31:0] c21;
wire[31:0] c22;
wire[31:0] c23;
wire[31:0] c24;
wire[31:0] c25;
wire[31:0] c26;
wire[31:0] c27;
wire[31:0] c28;
wire[31:0] c29;
wire[31:0] c30;
wire[31:0] c31;
wire[31:0] c32;
wire[31:0] c33;
wire[31:0] c34;
wire[31:0] c35;
wire[31:0] c36;
wire[31:0] c37;
wire[31:0] c38;
wire[31:0] c39;
wire[31:0] c40;
wire[31:0] c41;
wire[31:0] c42;
wire[31:0] c43;
wire[31:0] c44;
wire[31:0] c45;
wire[31:0] c46;
wire[31:0] c47;
wire[31:0] c48;
wire[31:0] c49;
wire[31:0] c50;
wire[31:0] c51;
wire[31:0] c52;
wire[31:0] c53;
wire[31:0] c54;
wire[31:0] c55;
wire[31:0] c56;
wire[31:0] c57;
wire[31:0] c58;
wire[31:0] c59;
wire[31:0] c60;
wire[31:0] c61;
wire[31:0] c62;
wire[31:0] c63;
wire[31:0] c64;
wire[31:0] c65;
wire[31:0] c66;
wire[31:0] c67;
wire[31:0] c68;
wire[31:0] c69;
wire[31:0] c70;
wire[31:0] c71;
wire[31:0] c72;
wire[31:0] c73;
wire[31:0] c74;
wire[31:0] c75;
wire[31:0] c76;
wire[31:0] c77;
wire[31:0] c78;
wire[31:0] c79;
wire[31:0] c80;
wire[31:0] d0;
wire[31:0] d1;
wire[31:0] d2;
wire[31:0] d3;
wire[31:0] d4;
wire[31:0] d5;
wire[31:0] d6;
wire[31:0] d7;
wire[31:0] d8;
wire[31:0] d9;
wire[31:0] d10;
wire[31:0] d11;
wire[31:0] d12;
wire[31:0] d13;
wire[31:0] d14;
wire[31:0] d15;
wire[31:0] d16;
wire[31:0] d17;
wire[31:0] d18;
wire[31:0] d19;
wire[31:0] d20;
wire[31:0] d21;
wire[31:0] d22;
wire[31:0] d23;
wire[31:0] d24;
wire[31:0] d25;
wire[31:0] d26;
wire[31:0] d27;
wire[31:0] d28;
wire[31:0] d29;
wire[31:0] d30;
wire[31:0] d31;
wire[31:0] d32;
wire[31:0] d33;
wire[31:0] d34;
wire[31:0] d35;
wire[31:0] d36;
wire[31:0] d37;
wire[31:0] d38;
wire[31:0] d39;
wire[31:0] d40;
wire[31:0] d41;
wire[31:0] d42;
wire[31:0] d43;
wire[31:0] d44;
wire[31:0] d45;
wire[31:0] d46;
wire[31:0] d47;
wire[31:0] d48;
wire[31:0] d49;
wire[31:0] d50;
wire[31:0] d51;
wire[31:0] d52;
wire[31:0] d53;
wire[31:0] d54;
wire[31:0] d55;
wire[31:0] d56;
wire[31:0] d57;
wire[31:0] d58;
wire[31:0] d59;
wire[31:0] d60;
wire[31:0] d61;
wire[31:0] d62;
wire[31:0] d63;
wire[31:0] d64;
wire[31:0] d65;
wire[31:0] d66;
wire[31:0] d67;
wire[31:0] d68;
wire[31:0] d69;
wire[31:0] d70;
wire[31:0] d71;
wire[31:0] d72;
wire[31:0] d73;
wire[31:0] d74;
wire[31:0] d75;
wire[31:0] d76;
wire[31:0] d77;
wire[31:0] d78;
wire[31:0] d79;
wire[31:0] d80;
wire[31:0] e0;
wire[31:0] e1;
wire[31:0] e2;
wire[31:0] e3;
wire[31:0] e4;
wire[31:0] e5;
wire[31:0] e6;
wire[31:0] e7;
wire[31:0] e8;
wire[31:0] e9;
wire[31:0] e10;
wire[31:0] e11;
wire[31:0] e12;
wire[31:0] e13;
wire[31:0] e14;
wire[31:0] e15;
wire[31:0] e16;
wire[31:0] e17;
wire[31:0] e18;
wire[31:0] e19;
wire[31:0] e20;
wire[31:0] e21;
wire[31:0] e22;
wire[31:0] e23;
wire[31:0] e24;
wire[31:0] e25;
wire[31:0] e26;
wire[31:0] e27;
wire[31:0] e28;
wire[31:0] e29;
wire[31:0] e30;
wire[31:0] e31;
wire[31:0] e32;
wire[31:0] e33;
wire[31:0] e34;
wire[31:0] e35;
wire[31:0] e36;
wire[31:0] e37;
wire[31:0] e38;
wire[31:0] e39;
wire[31:0] e40;
wire[31:0] e41;
wire[31:0] e42;
wire[31:0] e43;
wire[31:0] e44;
wire[31:0] e45;
wire[31:0] e46;
wire[31:0] e47;
wire[31:0] e48;
wire[31:0] e49;
wire[31:0] e50;
wire[31:0] e51;
wire[31:0] e52;
wire[31:0] e53;
wire[31:0] e54;
wire[31:0] e55;
wire[31:0] e56;
wire[31:0] e57;
wire[31:0] e58;
wire[31:0] e59;
wire[31:0] e60;
wire[31:0] e61;
wire[31:0] e62;
wire[31:0] e63;
wire[31:0] e64;
wire[31:0] e65;
wire[31:0] e66;
wire[31:0] e67;
wire[31:0] e68;
wire[31:0] e69;
wire[31:0] e70;
wire[31:0] e71;
wire[31:0] e72;
wire[31:0] e73;
wire[31:0] e74;
wire[31:0] e75;
wire[31:0] e76;
wire[31:0] e77;
wire[31:0] e78;
wire[31:0] e79;
wire[31:0] e80;
assign w0 = W[0];
assign w1 = W[1];
assign w2 = W[2];
assign w3 = W[3];
assign w4 = W[4];
assign w5 = W[5];
assign w6 = W[6];
assign w7 = W[7];
assign w8 = W[8];
assign w9 = W[9];
assign w10 = W[10];
assign w11 = W[11];
assign w12 = W[12];
assign w13 = W[13];
assign w14 = W[14];
assign w15 = W[15];
assign w16 = W[16];
assign w17 = W[17];
assign w18 = W[18];
assign w19 = W[19];
assign w20 = W[20];
assign w21 = W[21];
assign w22 = W[22];
assign w23 = W[23];
assign w24 = W[24];
assign w25 = W[25];
assign w26 = W[26];
assign w27 = W[27];
assign w28 = W[28];
assign w29 = W[29];
assign w30 = W[30];
assign w31 = W[31];
assign w32 = W[32];
assign w33 = W[33];
assign w34 = W[34];
assign w35 = W[35];
assign w36 = W[36];
assign w37 = W[37];
assign w38 = W[38];
assign w39 = W[39];
assign w40 = W[40];
assign w41 = W[41];
assign w42 = W[42];
assign w43 = W[43];
assign w44 = W[44];
assign w45 = W[45];
assign w46 = W[46];
assign w47 = W[47];
assign w48 = W[48];
assign w49 = W[49];
assign w50 = W[50];
assign w51 = W[51];
assign w52 = W[52];
assign w53 = W[53];
assign w54 = W[54];
assign w55 = W[55];
assign w56 = W[56];
assign w57 = W[57];
assign w58 = W[58];
assign w59 = W[59];
assign w60 = W[60];
assign w61 = W[61];
assign w62 = W[62];
assign w63 = W[63];
assign w64 = W[64];
assign w65 = W[65];
assign w66 = W[66];
assign w67 = W[67];
assign w68 = W[68];
assign w69 = W[69];
assign w70 = W[70];
assign w71 = W[71];
assign w72 = W[72];
assign w73 = W[73];
assign w74 = W[74];
assign w75 = W[75];
assign w76 = W[76];
assign w77 = W[77];
assign w78 = W[78];
assign w79 = W[79];
assign w80 = W[80];
assign a0 = A[0];
assign a1 = A[1];
assign a2 = A[2];
assign a3 = A[3];
assign a4 = A[4];
assign a5 = A[5];
assign a6 = A[6];
assign a7 = A[7];
assign a8 = A[8];
assign a9 = A[9];
assign a10 = A[10];
assign a11 = A[11];
assign a12 = A[12];
assign a13 = A[13];
assign a14 = A[14];
assign a15 = A[15];
assign a16 = A[16];
assign a17 = A[17];
assign a18 = A[18];
assign a19 = A[19];
assign a20 = A[20];
assign a21 = A[21];
assign a22 = A[22];
assign a23 = A[23];
assign a24 = A[24];
assign a25 = A[25];
assign a26 = A[26];
assign a27 = A[27];
assign a28 = A[28];
assign a29 = A[29];
assign a30 = A[30];
assign a31 = A[31];
assign a32 = A[32];
assign a33 = A[33];
assign a34 = A[34];
assign a35 = A[35];
assign a36 = A[36];
assign a37 = A[37];
assign a38 = A[38];
assign a39 = A[39];
assign a40 = A[40];
assign a41 = A[41];
assign a42 = A[42];
assign a43 = A[43];
assign a44 = A[44];
assign a45 = A[45];
assign a46 = A[46];
assign a47 = A[47];
assign a48 = A[48];
assign a49 = A[49];
assign a50 = A[50];
assign a51 = A[51];
assign a52 = A[52];
assign a53 = A[53];
assign a54 = A[54];
assign a55 = A[55];
assign a56 = A[56];
assign a57 = A[57];
assign a58 = A[58];
assign a59 = A[59];
assign a60 = A[60];
assign a61 = A[61];
assign a62 = A[62];
assign a63 = A[63];
assign a64 = A[64];
assign a65 = A[65];
assign a66 = A[66];
assign a67 = A[67];
assign a68 = A[68];
assign a69 = A[69];
assign a70 = A[70];
assign a71 = A[71];
assign a72 = A[72];
assign a73 = A[73];
assign a74 = A[74];
assign a75 = A[75];
assign a76 = A[76];
assign a77 = A[77];
assign a78 = A[78];
assign a79 = A[79];
assign a80 = A[80];
assign b0 = B[0];
assign b1 = B[1];
assign b2 = B[2];
assign b3 = B[3];
assign b4 = B[4];
assign b5 = B[5];
assign b6 = B[6];
assign b7 = B[7];
assign b8 = B[8];
assign b9 = B[9];
assign b10 = B[10];
assign b11 = B[11];
assign b12 = B[12];
assign b13 = B[13];
assign b14 = B[14];
assign b15 = B[15];
assign b16 = B[16];
assign b17 = B[17];
assign b18 = B[18];
assign b19 = B[19];
assign b20 = B[20];
assign b21 = B[21];
assign b22 = B[22];
assign b23 = B[23];
assign b24 = B[24];
assign b25 = B[25];
assign b26 = B[26];
assign b27 = B[27];
assign b28 = B[28];
assign b29 = B[29];
assign b30 = B[30];
assign b31 = B[31];
assign b32 = B[32];
assign b33 = B[33];
assign b34 = B[34];
assign b35 = B[35];
assign b36 = B[36];
assign b37 = B[37];
assign b38 = B[38];
assign b39 = B[39];
assign b40 = B[40];
assign b41 = B[41];
assign b42 = B[42];
assign b43 = B[43];
assign b44 = B[44];
assign b45 = B[45];
assign b46 = B[46];
assign b47 = B[47];
assign b48 = B[48];
assign b49 = B[49];
assign b50 = B[50];
assign b51 = B[51];
assign b52 = B[52];
assign b53 = B[53];
assign b54 = B[54];
assign b55 = B[55];
assign b56 = B[56];
assign b57 = B[57];
assign b58 = B[58];
assign b59 = B[59];
assign b60 = B[60];
assign b61 = B[61];
assign b62 = B[62];
assign b63 = B[63];
assign b64 = B[64];
assign b65 = B[65];
assign b66 = B[66];
assign b67 = B[67];
assign b68 = B[68];
assign b69 = B[69];
assign b70 = B[70];
assign b71 = B[71];
assign b72 = B[72];
assign b73 = B[73];
assign b74 = B[74];
assign b75 = B[75];
assign b76 = B[76];
assign b77 = B[77];
assign b78 = B[78];
assign b79 = B[79];
assign b80 = B[80];
assign c0 = C[0];
assign c1 = C[1];
assign c2 = C[2];
assign c3 = C[3];
assign c4 = C[4];
assign c5 = C[5];
assign c6 = C[6];
assign c7 = C[7];
assign c8 = C[8];
assign c9 = C[9];
assign c10 = C[10];
assign c11 = C[11];
assign c12 = C[12];
assign c13 = C[13];
assign c14 = C[14];
assign c15 = C[15];
assign c16 = C[16];
assign c17 = C[17];
assign c18 = C[18];
assign c19 = C[19];
assign c20 = C[20];
assign c21 = C[21];
assign c22 = C[22];
assign c23 = C[23];
assign c24 = C[24];
assign c25 = C[25];
assign c26 = C[26];
assign c27 = C[27];
assign c28 = C[28];
assign c29 = C[29];
assign c30 = C[30];
assign c31 = C[31];
assign c32 = C[32];
assign c33 = C[33];
assign c34 = C[34];
assign c35 = C[35];
assign c36 = C[36];
assign c37 = C[37];
assign c38 = C[38];
assign c39 = C[39];
assign c40 = C[40];
assign c41 = C[41];
assign c42 = C[42];
assign c43 = C[43];
assign c44 = C[44];
assign c45 = C[45];
assign c46 = C[46];
assign c47 = C[47];
assign c48 = C[48];
assign c49 = C[49];
assign c50 = C[50];
assign c51 = C[51];
assign c52 = C[52];
assign c53 = C[53];
assign c54 = C[54];
assign c55 = C[55];
assign c56 = C[56];
assign c57 = C[57];
assign c58 = C[58];
assign c59 = C[59];
assign c60 = C[60];
assign c61 = C[61];
assign c62 = C[62];
assign c63 = C[63];
assign c64 = C[64];
assign c65 = C[65];
assign c66 = C[66];
assign c67 = C[67];
assign c68 = C[68];
assign c69 = C[69];
assign c70 = C[70];
assign c71 = C[71];
assign c72 = C[72];
assign c73 = C[73];
assign c74 = C[74];
assign c75 = C[75];
assign c76 = C[76];
assign c77 = C[77];
assign c78 = C[78];
assign c79 = C[79];
assign c80 = C[80];
assign d0 = D[0];
assign d1 = D[1];
assign d2 = D[2];
assign d3 = D[3];
assign d4 = D[4];
assign d5 = D[5];
assign d6 = D[6];
assign d7 = D[7];
assign d8 = D[8];
assign d9 = D[9];
assign d10 = D[10];
assign d11 = D[11];
assign d12 = D[12];
assign d13 = D[13];
assign d14 = D[14];
assign d15 = D[15];
assign d16 = D[16];
assign d17 = D[17];
assign d18 = D[18];
assign d19 = D[19];
assign d20 = D[20];
assign d21 = D[21];
assign d22 = D[22];
assign d23 = D[23];
assign d24 = D[24];
assign d25 = D[25];
assign d26 = D[26];
assign d27 = D[27];
assign d28 = D[28];
assign d29 = D[29];
assign d30 = D[30];
assign d31 = D[31];
assign d32 = D[32];
assign d33 = D[33];
assign d34 = D[34];
assign d35 = D[35];
assign d36 = D[36];
assign d37 = D[37];
assign d38 = D[38];
assign d39 = D[39];
assign d40 = D[40];
assign d41 = D[41];
assign d42 = D[42];
assign d43 = D[43];
assign d44 = D[44];
assign d45 = D[45];
assign d46 = D[46];
assign d47 = D[47];
assign d48 = D[48];
assign d49 = D[49];
assign d50 = D[50];
assign d51 = D[51];
assign d52 = D[52];
assign d53 = D[53];
assign d54 = D[54];
assign d55 = D[55];
assign d56 = D[56];
assign d57 = D[57];
assign d58 = D[58];
assign d59 = D[59];
assign d60 = D[60];
assign d61 = D[61];
assign d62 = D[62];
assign d63 = D[63];
assign d64 = D[64];
assign d65 = D[65];
assign d66 = D[66];
assign d67 = D[67];
assign d68 = D[68];
assign d69 = D[69];
assign d70 = D[70];
assign d71 = D[71];
assign d72 = D[72];
assign d73 = D[73];
assign d74 = D[74];
assign d75 = D[75];
assign d76 = D[76];
assign d77 = D[77];
assign d78 = D[78];
assign d79 = D[79];
assign d80 = D[80];
assign e0 = E[0];
assign e1 = E[1];
assign e2 = E[2];
assign e3 = E[3];
assign e4 = E[4];
assign e5 = E[5];
assign e6 = E[6];
assign e7 = E[7];
assign e8 = E[8];
assign e9 = E[9];
assign e10 = E[10];
assign e11 = E[11];
assign e12 = E[12];
assign e13 = E[13];
assign e14 = E[14];
assign e15 = E[15];
assign e16 = E[16];
assign e17 = E[17];
assign e18 = E[18];
assign e19 = E[19];
assign e20 = E[20];
assign e21 = E[21];
assign e22 = E[22];
assign e23 = E[23];
assign e24 = E[24];
assign e25 = E[25];
assign e26 = E[26];
assign e27 = E[27];
assign e28 = E[28];
assign e29 = E[29];
assign e30 = E[30];
assign e31 = E[31];
assign e32 = E[32];
assign e33 = E[33];
assign e34 = E[34];
assign e35 = E[35];
assign e36 = E[36];
assign e37 = E[37];
assign e38 = E[38];
assign e39 = E[39];
assign e40 = E[40];
assign e41 = E[41];
assign e42 = E[42];
assign e43 = E[43];
assign e44 = E[44];
assign e45 = E[45];
assign e46 = E[46];
assign e47 = E[47];
assign e48 = E[48];
assign e49 = E[49];
assign e50 = E[50];
assign e51 = E[51];
assign e52 = E[52];
assign e53 = E[53];
assign e54 = E[54];
assign e55 = E[55];
assign e56 = E[56];
assign e57 = E[57];
assign e58 = E[58];
assign e59 = E[59];
assign e60 = E[60];
assign e61 = E[61];
assign e62 = E[62];
assign e63 = E[63];
assign e64 = E[64];
assign e65 = E[65];
assign e66 = E[66];
assign e67 = E[67];
assign e68 = E[68];
assign e69 = E[69];
assign e70 = E[70];
assign e71 = E[71];
assign e72 = E[72];
assign e73 = E[73];
assign e74 = E[74];
assign e75 = E[75];
assign e76 = E[76];
assign e77 = E[77];
assign e78 = E[78];
assign e79 = E[79];
assign e80 = E[80];


    integer i;
    always @(*) begin
        sha_pad[63:0] <= 64'd32;
        sha_pad[511:480] <= sha1_i;
        sha_pad[478:64] <= 415'd0;
        sha_pad[479] <= 1;
        A[0] <= 32'h67452301;
        B[0] <= 32'hEFCDAB89;
        C[0] <= 32'h98BADCFE;
        D[0] <= 32'h10325476;
        E[0] <= 32'hC3D2E1F0;
        W[1] <= sha_pad[511:480];
        W[2] <= sha_pad[479:448];
        W[3] <= sha_pad[447:416];
        W[4] <= sha_pad[415:384];
        W[5] <= sha_pad[383:352];
        W[6] <= sha_pad[351:320];
        W[7] <= sha_pad[319:288];
        W[8] <= sha_pad[287:256];
        W[9] <= sha_pad[255:224];
        W[10] <= sha_pad[223:192];
        W[11] <= sha_pad[191:160];
        W[12] <= sha_pad[159:128];
        W[13] <= sha_pad[127:96];
        W[14] <= sha_pad[95:64];
        W[15] <= sha_pad[63:32];
        W[16] <= sha_pad[31:0];
        for (i = 1; i<=16; i=i+1) begin
            A[i] <= ((A[i-1]<<5)|(A[i-1]>>(32-5))) + ((B[i-1]&C[i-1])|((~B[i-1]) & D[i-1])) + (E[i-1]) +W[i] + 32'h5A827999;
            E[i] <= D[i-1];
            D[i] <= C[i-1];
            C[i] <= ((B[i-1]<<30)|(B[i-1]>>2));
            B[i] <= A[i-1];
        end

        for (i = 17; i<=20; i=i+1) begin
            W[i] <= ((W[i-3]^W[i-8]^W[i-14]^W[i-16])<<1)|((W[i-3]^W[i-8]^W[i-14]^W[i-16])>>31);
            A[i] <= ((A[i-1]<<5)|(A[i-1]>>(32-5))) + ((B[i-1]&C[i-1])|((~B[i-1]) & D[i-1])) + (E[i-1]) +W[i] + 32'h5A827999;
            E[i] <= D[i-1];
            D[i] <= C[i-1];
            C[i] <= ((B[i-1]<<30)|(B[i-1]>>2));
            B[i] <= A[i-1];
        end
        for (i = 21; i<=40; i=i+1) begin
            W[i] <= ((W[i-3]^W[i-8]^W[i-14]^W[i-16])<<1)|((W[i-3]^W[i-8]^W[i-14]^W[i-16])>>31);
            A[i] <= ((A[i-1]<<5)|(A[i-1]>>(32-5))) + (B[i-1]^C[i-1]^D[i-1]) + (E[i-1]) +W[i] + 32'h6ED9EBA1;
            E[i] <= D[i-1];
            D[i] <= C[i-1];
            C[i] <= ((B[i-1]<<30)|(B[i-1]>>2));
            B[i] <= A[i-1];
        end

        for (i = 41; i<=60; i=i+1) begin
            W[i] <= ((W[i-3]^W[i-8]^W[i-14]^W[i-16])<<1)|((W[i-3]^W[i-8]^W[i-14]^W[i-16])>>31);
            A[i] <= ((A[i-1]<<5)|(A[i-1]>>(32-5))) + ((B[i-1]&C[i-1])|(B[i-1]&D[i-1])|(C[i-1]&D[i-1]))+ (E[i-1]) +W[i] + 32'h8F1BBCDC;
            E[i] <= D[i-1];
            D[i] <= C[i-1];
            C[i] <= ((B[i-1]<<30)|(B[i-1]>>2));
            B[i] <= A[i-1];
        end

        for (i = 61; i<=80; i=i+1) begin
            W[i] <= ((W[i-3]^W[i-8]^W[i-14]^W[i-16])<<1)|((W[i-3]^W[i-8]^W[i-14]^W[i-16])>>31);
            A[i] <= ((A[i-1]<<5)|(A[i-1]>>(32-5))) + (B[i-1]^C[i-1]^D[i-1]) + (E[i-1]) +W[i] + 32'hCA62C1D6;
            E[i] <= D[i-1];
            D[i] <= C[i-1];
            C[i] <= ((B[i-1]<<30)|(B[i-1]>>2));
            B[i] <= A[i-1];
        end
        // sha1_o[159:128] <= A[0] + A[80];
        // sha1_o[127:96] <= B[0] + B[80];
        // sha1_o[95:64] <= C[0] + C[80];
        // sha1_o[63:32] <= D[0] + D[80];
        // sha1_o[32:0] <= E[0] + E[80];
    end


    // for (i = 21; i<=40; i=i+1) begin
    //     assign W[i] = ((W[i-3]^W[i-8]^W[i-14]^W[i-16])<<1)|((W[i-3]^W[i-8]^W[i-14]^W[i-16])>>31);
    //     assign A[i] = ((A[i-1]<<5)|(A[i-1]>>(32-5))) + (B[i-1]&C[i-1])|(B[i-1]&D[i-1])|(C[i-1]&D[i-1]) + (E[i-1]) +W[i] + 32'h6ED9EBA1;
    //     assign E[i] = D[i-1];
    //     assign D[i] = C[i-1];
    //     assign C[i] = ((B[i-1]<<30)|(B[i-1]>>2));
    //     assign B[i] = A[i-1];
    // end

    // for (i = 41; i<=60; i=i+1) begin
    //     assign W[i] = ((W[i-3]^W[i-8]^W[i-14]^W[i-16])<<1)|((W[i-3]^W[i-8]^W[i-14]^W[i-16])>>31);
    //     assign A[i] = ((A[i-1]<<5)|(A[i-1]>>(32-5))) +(B[i-1]^C[i-1]^D[i-1])+ (E[i-1]) +W[i] + 32'h8F1BBCDC;
    //     assign E[i] = D[i-1];
    //     assign D[i] = C[i-1];
    //     assign C[i] = ((B[i-1]<<30)|(B[i-1]>>2));
    //     assign B[i] = A[i-1];
    // end

    // for (i = 61; i<=80; i=i+1) begin
    //     assign W[i] = ((W[i-3]^W[i-8]^W[i-14]^W[i-16])<<1)|((W[i-3]^W[i-8]^W[i-14]^W[i-16])>>31);
    //     assign A[i] = ((A[i-1]<<5)|(A[i-1]>>(32-5))) + (B[i-1]&C[i-1])|(B[i-1]&D[i-1])|(C[i-1]&D[i-1]) + (E[i-1]) +W[i] + 32'hCA62C1D6;
    //     assign E[i] = D[i-1];
    //     assign D[i] = C[i-1];
    //     assign C[i] = ((B[i-1]<<30)|(B[i-1]>>2));
    //     assign B[i] = A[i-1];
    // end

    assign sha1_o[159:128] = A[0] + A[80];
    assign sha1_o[127:96] = B[0] + B[80];
    assign sha1_o[95:64] = C[0] + C[80];
    assign sha1_o[63:32] = D[0] + D[80];
    assign sha1_o[31:0] = E[0] + E[80];

endmodule


// module fun1(

//     input wire B[31:0],
//     input wire C[31:0],
//     input wire D[31:0],
//     output wire O[31:0]
//     );

//     assign O = (B & C) | ((~B) & D);

// endmodule

// module fun2(

//     input wire B[31:0],
//     input wire C[31:0],
//     input wire D[31:0],
//     output wire O[31:0]
//     );

//     assign O = B ^ C ^ D;

// endmodule

// module fun3(

//     input wire B[31:0],
//     input wire C[31:0],
//     input wire D[31:0],
//     output wire O[31:0]
//     );

//     assign O = (B & C) | (B & D) | (C & D);

// endmodule

// module fun4(

//     input wire B[31:0],
//     input wire C[31:0],
//     input wire D[31:0],
//     output wire O[31:0]
//     );

//     assign O = (B & C) | (B & D) | (C & D);

// endmodule